module RnG(
input wire [1:0] state,
input wire clk,
output wire [4:0] RnG
);
	reg [4:0] counter;        
	reg [4:0] RnG_reg;
	reg [4:0] RnG_reg2;



	
	
endmodule